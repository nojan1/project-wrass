module top (

)  
